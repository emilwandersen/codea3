module DataMemory(
  input         clock,
  input  [15:0] io_address,
  output [31:0] io_dataRead,
  input         io_writeEnable,
  input  [31:0] io_dataWrite,
  input         io_testerEnable,
  input  [15:0] io_testerAddress,
  output [31:0] io_testerDataRead,
  input         io_testerWriteEnable,
  input  [31:0] io_testerDataWrite
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
  reg [31:0] memory [0:65535]; // @[DataMemory.scala 18:20]
  wire [31:0] memory__T_data; // @[DataMemory.scala 18:20]
  wire [15:0] memory__T_addr; // @[DataMemory.scala 18:20]
  wire [31:0] memory__T_2_data; // @[DataMemory.scala 18:20]
  wire [15:0] memory__T_2_addr; // @[DataMemory.scala 18:20]
  wire [31:0] memory__T_1_data; // @[DataMemory.scala 18:20]
  wire [15:0] memory__T_1_addr; // @[DataMemory.scala 18:20]
  wire  memory__T_1_mask; // @[DataMemory.scala 18:20]
  wire  memory__T_1_en; // @[DataMemory.scala 18:20]
  wire [31:0] memory__T_3_data; // @[DataMemory.scala 18:20]
  wire [15:0] memory__T_3_addr; // @[DataMemory.scala 18:20]
  wire  memory__T_3_mask; // @[DataMemory.scala 18:20]
  wire  memory__T_3_en; // @[DataMemory.scala 18:20]
  wire [31:0] _GEN_5 = io_testerWriteEnable ? io_testerDataWrite : memory__T_data; // @[DataMemory.scala 27:32]
  wire [31:0] _GEN_11 = io_writeEnable ? io_dataWrite : memory__T_2_data; // @[DataMemory.scala 37:26]
  assign memory__T_addr = io_testerAddress;
  assign memory__T_data = memory[memory__T_addr]; // @[DataMemory.scala 18:20]
  assign memory__T_2_addr = io_address;
  assign memory__T_2_data = memory[memory__T_2_addr]; // @[DataMemory.scala 18:20]
  assign memory__T_1_data = io_testerDataWrite;
  assign memory__T_1_addr = io_testerAddress;
  assign memory__T_1_mask = 1'h1;
  assign memory__T_1_en = io_testerEnable & io_testerWriteEnable;
  assign memory__T_3_data = io_dataWrite;
  assign memory__T_3_addr = io_address;
  assign memory__T_3_mask = 1'h1;
  assign memory__T_3_en = io_testerEnable ? 1'h0 : io_writeEnable;
  assign io_dataRead = io_testerEnable ? 32'h0 : _GEN_11; // @[DataMemory.scala 26:17 DataMemory.scala 34:17 DataMemory.scala 40:19]
  assign io_testerDataRead = io_testerEnable ? _GEN_5 : 32'h0; // @[DataMemory.scala 24:23 DataMemory.scala 30:25 DataMemory.scala 36:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 65536; initvar = initvar+1)
    memory[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(memory__T_1_en & memory__T_1_mask) begin
      memory[memory__T_1_addr] <= memory__T_1_data; // @[DataMemory.scala 18:20]
    end
    if(memory__T_3_en & memory__T_3_mask) begin
      memory[memory__T_3_addr] <= memory__T_3_data; // @[DataMemory.scala 18:20]
    end
  end
endmodule
module Accelerator(
  input         clock,
  input         reset,
  input         io_start,
  output        io_done,
  output [15:0] io_address,
  input  [31:0] io_dataRead,
  output        io_writeEnable,
  output [31:0] io_dataWrite
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] x; // @[Accelerator.scala 26:18]
  reg [15:0] y; // @[Accelerator.scala 27:18]
  reg [31:0] in; // @[Accelerator.scala 28:19]
  reg [31:0] op; // @[Accelerator.scala 29:19]
  reg [31:0] value; // @[Accelerator.scala 30:21]
  reg [31:0] left; // @[Accelerator.scala 31:21]
  reg [31:0] right; // @[Accelerator.scala 32:21]
  reg [31:0] up; // @[Accelerator.scala 33:19]
  reg [31:0] down; // @[Accelerator.scala 34:21]
  reg [3:0] stateReg; // @[Accelerator.scala 40:25]
  wire  _T = 4'h1 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_1 = 4'h0 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_2 = 4'h2 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_3 = x < 16'h14; // @[Accelerator.scala 64:13]
  wire  _T_4 = 4'h3 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_5 = y < 16'h14; // @[Accelerator.scala 74:13]
  wire  _T_6 = x == 16'h0; // @[Accelerator.scala 76:15]
  wire  _T_7 = y == 16'h0; // @[Accelerator.scala 76:23]
  wire  _T_8 = _T_6 | _T_7; // @[Accelerator.scala 76:21]
  wire  _T_9 = x == 16'h13; // @[Accelerator.scala 76:31]
  wire  _T_10 = _T_8 | _T_9; // @[Accelerator.scala 76:29]
  wire  _T_11 = y == 16'h13; // @[Accelerator.scala 76:40]
  wire  _T_12 = _T_10 | _T_11; // @[Accelerator.scala 76:38]
  wire [15:0] _T_14 = x + 16'h1; // @[Accelerator.scala 85:14]
  wire  _T_15 = 4'h4 == stateReg; // @[Conditional.scala 37:30]
  wire [15:0] _T_17 = y + 16'h1; // @[Accelerator.scala 94:11]
  wire [31:0] _T_19 = op + 32'h1; // @[Accelerator.scala 95:13]
  wire [31:0] _T_21 = in + 32'h1; // @[Accelerator.scala 96:13]
  wire  _T_22 = 4'h5 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_29 = 4'h6 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_30 = 4'h7 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_31 = value == 32'h0; // @[Accelerator.scala 116:17]
  wire [31:0] _T_33 = in - 32'h1; // @[Accelerator.scala 119:23]
  wire [31:0] _GEN_7 = _T_31 ? 32'h0 : _T_33; // @[Accelerator.scala 116:24]
  wire  _T_34 = 4'h8 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_35 = left == 32'h0; // @[Accelerator.scala 125:16]
  wire [31:0] _GEN_10 = _T_35 ? 32'h0 : _T_21; // @[Accelerator.scala 125:23]
  wire  _T_38 = 4'h9 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_39 = right == 32'h0; // @[Accelerator.scala 134:18]
  wire [31:0] _T_41 = in - 32'h14; // @[Accelerator.scala 137:26]
  wire [31:0] _GEN_13 = _T_39 ? 32'h0 : _T_41; // @[Accelerator.scala 134:27]
  wire  _T_42 = 4'ha == stateReg; // @[Conditional.scala 37:30]
  wire  _T_43 = up == 32'h0; // @[Accelerator.scala 144:15]
  wire [31:0] _T_45 = in + 32'h14; // @[Accelerator.scala 147:26]
  wire [31:0] _GEN_16 = _T_43 ? 32'h0 : _T_45; // @[Accelerator.scala 144:24]
  wire  _T_46 = 4'hb == stateReg; // @[Conditional.scala 37:30]
  wire  _T_47 = down == 32'h0; // @[Accelerator.scala 153:16]
  wire [31:0] _GEN_21 = _T_42 ? _GEN_16 : 32'h0; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_24 = _T_38 ? _GEN_13 : _GEN_21; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_28 = _T_34 ? _GEN_10 : _GEN_24; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_33 = _T_30 ? _GEN_7 : _GEN_28; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_38 = _T_29 ? in : _GEN_33; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_45 = _T_22 ? op : _GEN_38; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_47 = _T_22 ? 8'hff : 8'h0; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_57 = _T_15 ? op : _GEN_45; // @[Conditional.scala 39:67]
  wire  _GEN_58 = _T_15 | _T_22; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_59 = _T_15 ? 8'h0 : _GEN_47; // @[Conditional.scala 39:67]
  wire  _GEN_69 = _T_4 ? 1'h0 : _GEN_58; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_72 = _T_4 ? 32'h0 : _GEN_57; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_73 = _T_4 ? 8'h0 : _GEN_59; // @[Conditional.scala 39:67]
  wire  _GEN_84 = _T_2 ? 1'h0 : _GEN_69; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_86 = _T_2 ? 32'h0 : _GEN_72; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_87 = _T_2 ? 8'h0 : _GEN_73; // @[Conditional.scala 39:67]
  wire  _GEN_100 = _T_1 ? 1'h0 : _GEN_84; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_101 = _T_1 ? 32'h0 : _GEN_86; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_102 = _T_1 ? 8'h0 : _GEN_87; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_115 = _T ? 32'h0 : _GEN_101; // @[Conditional.scala 40:58]
  wire [7:0] _GEN_116 = _T ? 8'h0 : _GEN_102; // @[Conditional.scala 40:58]
  assign io_done = 4'h1 == stateReg; // @[Accelerator.scala 21:10 Accelerator.scala 50:14]
  assign io_address = _GEN_115[15:0]; // @[Accelerator.scala 22:13 Accelerator.scala 91:17 Accelerator.scala 101:18 Accelerator.scala 111:17 Accelerator.scala 119:19 Accelerator.scala 128:19 Accelerator.scala 137:20 Accelerator.scala 147:20]
  assign io_writeEnable = _T ? 1'h0 : _GEN_100; // @[Accelerator.scala 23:17 Accelerator.scala 73:21 Accelerator.scala 92:21 Accelerator.scala 102:22]
  assign io_dataWrite = {{24'd0}, _GEN_116}; // @[Accelerator.scala 24:15 Accelerator.scala 93:19 Accelerator.scala 103:20]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  x = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  y = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  in = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  op = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  value = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  left = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  right = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  up = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  down = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  stateReg = _RAND_9[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      x <= 16'h0;
    end else if (!(_T)) begin
      if (_T_1) begin
        x <= 16'h0;
      end else if (!(_T_2)) begin
        if (_T_4) begin
          if (!(_T_5)) begin
            x <= _T_14;
          end
        end
      end
    end
    if (reset) begin
      y <= 16'h0;
    end else if (!(_T)) begin
      if (_T_1) begin
        y <= 16'h0;
      end else if (_T_2) begin
        if (_T_3) begin
          y <= 16'h0;
        end
      end else if (!(_T_4)) begin
        if (_T_15) begin
          y <= _T_17;
        end else if (_T_22) begin
          y <= _T_17;
        end
      end
    end
    if (reset) begin
      in <= 32'h0;
    end else if (!(_T)) begin
      if (_T_1) begin
        in <= 32'h0;
      end else if (!(_T_2)) begin
        if (!(_T_4)) begin
          if (_T_15) begin
            in <= _T_21;
          end else if (_T_22) begin
            in <= _T_21;
          end
        end
      end
    end
    if (reset) begin
      op <= 32'h190;
    end else if (!(_T)) begin
      if (_T_1) begin
        op <= 32'h190;
      end else if (!(_T_2)) begin
        if (!(_T_4)) begin
          if (_T_15) begin
            op <= _T_19;
          end else if (_T_22) begin
            op <= _T_19;
          end
        end
      end
    end
    if (reset) begin
      value <= 32'h0;
    end else if (!(_T)) begin
      if (!(_T_1)) begin
        if (!(_T_2)) begin
          if (!(_T_4)) begin
            if (!(_T_15)) begin
              if (!(_T_22)) begin
                if (_T_29) begin
                  value <= io_dataRead;
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      left <= 32'h0;
    end else if (!(_T)) begin
      if (!(_T_1)) begin
        if (!(_T_2)) begin
          if (!(_T_4)) begin
            if (!(_T_15)) begin
              if (!(_T_22)) begin
                if (!(_T_29)) begin
                  if (_T_30) begin
                    if (!(_T_31)) begin
                      left <= io_dataRead;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      right <= 32'h0;
    end else if (!(_T)) begin
      if (!(_T_1)) begin
        if (!(_T_2)) begin
          if (!(_T_4)) begin
            if (!(_T_15)) begin
              if (!(_T_22)) begin
                if (!(_T_29)) begin
                  if (!(_T_30)) begin
                    if (_T_34) begin
                      if (!(_T_35)) begin
                        right <= io_dataRead;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      up <= 32'h0;
    end else if (!(_T)) begin
      if (!(_T_1)) begin
        if (!(_T_2)) begin
          if (!(_T_4)) begin
            if (!(_T_15)) begin
              if (!(_T_22)) begin
                if (!(_T_29)) begin
                  if (!(_T_30)) begin
                    if (!(_T_34)) begin
                      if (_T_38) begin
                        if (!(_T_39)) begin
                          up <= io_dataRead;
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      down <= 32'h0;
    end else if (!(_T)) begin
      if (!(_T_1)) begin
        if (!(_T_2)) begin
          if (!(_T_4)) begin
            if (!(_T_15)) begin
              if (!(_T_22)) begin
                if (!(_T_29)) begin
                  if (!(_T_30)) begin
                    if (!(_T_34)) begin
                      if (!(_T_38)) begin
                        if (_T_42) begin
                          if (!(_T_43)) begin
                            down <= io_dataRead;
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      stateReg <= 4'h0;
    end else if (!(_T)) begin
      if (_T_1) begin
        if (io_start) begin
          stateReg <= 4'h2;
        end
      end else if (_T_2) begin
        if (_T_3) begin
          stateReg <= 4'h3;
        end else begin
          stateReg <= 4'h1;
        end
      end else if (_T_4) begin
        if (_T_5) begin
          if (_T_12) begin
            stateReg <= 4'h4;
          end else begin
            stateReg <= 4'h6;
          end
        end else begin
          stateReg <= 4'h2;
        end
      end else if (_T_15) begin
        stateReg <= 4'h3;
      end else if (_T_22) begin
        stateReg <= 4'h3;
      end else if (_T_29) begin
        stateReg <= 4'h7;
      end else if (_T_30) begin
        if (_T_31) begin
          stateReg <= 4'h4;
        end else begin
          stateReg <= 4'h8;
        end
      end else if (_T_34) begin
        if (_T_35) begin
          stateReg <= 4'h4;
        end else begin
          stateReg <= 4'h9;
        end
      end else if (_T_38) begin
        if (_T_39) begin
          stateReg <= 4'h4;
        end else begin
          stateReg <= 4'ha;
        end
      end else if (_T_42) begin
        if (_T_43) begin
          stateReg <= 4'h4;
        end else begin
          stateReg <= 4'hb;
        end
      end else if (_T_46) begin
        if (_T_47) begin
          stateReg <= 4'h4;
        end else begin
          stateReg <= 4'h5;
        end
      end
    end
  end
endmodule
module SystemTop(
  input         clock,
  input         reset,
  output        io_done,
  input         io_start,
  input         io_testerDataMemEnable,
  input  [15:0] io_testerDataMemAddress,
  output [31:0] io_testerDataMemDataRead,
  input         io_testerDataMemWriteEnable,
  input  [31:0] io_testerDataMemDataWrite
);
  wire  dataMemory_clock; // @[SystemTop.scala 18:26]
  wire [15:0] dataMemory_io_address; // @[SystemTop.scala 18:26]
  wire [31:0] dataMemory_io_dataRead; // @[SystemTop.scala 18:26]
  wire  dataMemory_io_writeEnable; // @[SystemTop.scala 18:26]
  wire [31:0] dataMemory_io_dataWrite; // @[SystemTop.scala 18:26]
  wire  dataMemory_io_testerEnable; // @[SystemTop.scala 18:26]
  wire [15:0] dataMemory_io_testerAddress; // @[SystemTop.scala 18:26]
  wire [31:0] dataMemory_io_testerDataRead; // @[SystemTop.scala 18:26]
  wire  dataMemory_io_testerWriteEnable; // @[SystemTop.scala 18:26]
  wire [31:0] dataMemory_io_testerDataWrite; // @[SystemTop.scala 18:26]
  wire  accelerator_clock; // @[SystemTop.scala 19:27]
  wire  accelerator_reset; // @[SystemTop.scala 19:27]
  wire  accelerator_io_start; // @[SystemTop.scala 19:27]
  wire  accelerator_io_done; // @[SystemTop.scala 19:27]
  wire [15:0] accelerator_io_address; // @[SystemTop.scala 19:27]
  wire [31:0] accelerator_io_dataRead; // @[SystemTop.scala 19:27]
  wire  accelerator_io_writeEnable; // @[SystemTop.scala 19:27]
  wire [31:0] accelerator_io_dataWrite; // @[SystemTop.scala 19:27]
  DataMemory dataMemory ( // @[SystemTop.scala 18:26]
    .clock(dataMemory_clock),
    .io_address(dataMemory_io_address),
    .io_dataRead(dataMemory_io_dataRead),
    .io_writeEnable(dataMemory_io_writeEnable),
    .io_dataWrite(dataMemory_io_dataWrite),
    .io_testerEnable(dataMemory_io_testerEnable),
    .io_testerAddress(dataMemory_io_testerAddress),
    .io_testerDataRead(dataMemory_io_testerDataRead),
    .io_testerWriteEnable(dataMemory_io_testerWriteEnable),
    .io_testerDataWrite(dataMemory_io_testerDataWrite)
  );
  Accelerator accelerator ( // @[SystemTop.scala 19:27]
    .clock(accelerator_clock),
    .reset(accelerator_reset),
    .io_start(accelerator_io_start),
    .io_done(accelerator_io_done),
    .io_address(accelerator_io_address),
    .io_dataRead(accelerator_io_dataRead),
    .io_writeEnable(accelerator_io_writeEnable),
    .io_dataWrite(accelerator_io_dataWrite)
  );
  assign io_done = accelerator_io_done; // @[SystemTop.scala 23:11]
  assign io_testerDataMemDataRead = dataMemory_io_testerDataRead; // @[SystemTop.scala 34:28]
  assign dataMemory_clock = clock;
  assign dataMemory_io_address = accelerator_io_address; // @[SystemTop.scala 28:25]
  assign dataMemory_io_writeEnable = accelerator_io_writeEnable; // @[SystemTop.scala 30:29]
  assign dataMemory_io_dataWrite = accelerator_io_dataWrite; // @[SystemTop.scala 29:27]
  assign dataMemory_io_testerEnable = io_testerDataMemEnable; // @[SystemTop.scala 36:30]
  assign dataMemory_io_testerAddress = io_testerDataMemAddress; // @[SystemTop.scala 33:31]
  assign dataMemory_io_testerWriteEnable = io_testerDataMemWriteEnable; // @[SystemTop.scala 37:35]
  assign dataMemory_io_testerDataWrite = io_testerDataMemDataWrite; // @[SystemTop.scala 35:33]
  assign accelerator_clock = clock;
  assign accelerator_reset = reset;
  assign accelerator_io_start = io_start; // @[SystemTop.scala 24:24]
  assign accelerator_io_dataRead = dataMemory_io_dataRead; // @[SystemTop.scala 27:27]
endmodule
